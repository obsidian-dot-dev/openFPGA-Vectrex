library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity compressor_lut is
port (
	data      : in  std_logic_vector(7 downto 0);
	data_comp : out std_logic_vector(5 downto 0)
);
end entity;

architecture prom of compressor_lut is
	type rom is array(0 to  255) of std_logic_vector(5 downto 0);
	signal rom_data: rom := (
	"000000","000000","000000","000000","000000","000000","000000","000001",
	"000001","000001","000001","000001","000001","000001","000001","000001",
	"000010","000010","000010","000010","000010","000010","000010","000011",
	"000011","000011","000011","000011","000011","000011","000100","000100",
	"000100","000100","000100","000100","000101","000101","000101","000101",
	"000101","000110","000110","000110","000110","000110","000110","000111",
	"000111","000111","000111","000111","001000","001000","001000","001000",
	"001000","001001","001001","001001","001001","001001","001010","001010",
	"001010","001010","001010","001011","001011","001011","001011","001011",
	"001100","001100","001100","001100","001101","001101","001101","001101",
	"001101","001110","001110","001110","001110","001111","001111","001111",
	"001111","001111","010000","010000","010000","010000","010001","010001",
	"010001","010001","010010","010010","010010","010010","010011","010011",
	"010011","010011","010100","010100","010100","010100","010101","010101",
	"010101","010101","010110","010110","010110","010110","010111","010111",
	"010111","010111","011000","011000","011000","011000","011001","011001",
	"011001","011001","011010","011010","011010","011010","011011","011011",
	"011011","011100","011100","011100","011100","011101","011101","011101",
	"011101","011110","011110","011110","011111","011111","011111","011111",
	"100000","100000","100000","100000","100001","100001","100001","100010",
	"100010","100010","100010","100011","100011","100011","100100","100100",
	"100100","100100","100101","100101","100101","100110","100110","100110",
	"100110","100111","100111","100111","101000","101000","101000","101000",
	"101001","101001","101001","101010","101010","101010","101011","101011",
	"101011","101011","101100","101100","101100","101101","101101","101101",
	"101110","101110","101110","101110","101111","101111","101111","110000",
	"110000","110000","110001","110001","110001","110010","110010","110010",
	"110010","110011","110011","110011","110100","110100","110100","110101",
	"110101","110101","110110","110110","110110","110111","110111","110111",
	"111000","111000","111000","111000","111001","111001","111001","111010",
	"111010","111010","111011","111011","111011","111100","111100","111100",
	"111101","111101","111101","111110","111110","111110","111111","111111"
  );
begin
data_comp <= rom_data(to_integer(unsigned(data)));
end architecture;
